module notm (
    input wire A, B,
    output wire C
    );
    assign C = A & B ;
endmodule